module hello;
initial begin
$display("Hello world");
end
endmodule
